128 720 660 47 978 360 222 299 842 831 757 550 429 53 533 306 767 30 767 230 555 389 858 724 953 998 850 714 49 395 883 860 508 529 884 800 809 430 33 613 269 522 295 307 105 764 221 667 965 93 239 992 265 517 788 526 697 289 652 645 837 397 528 732 578 835 194 511 914 818 167 984 485 268 382 265 44 380 206 915 62 470 897 542 902 374 443 365 447 434 297 749 217 908 295 664 67 359 772 37 313 886 738 431 348 501 563 282 164 273 502 60 477 180 602 468 45 656 324 880 444 947 380 71 697 982 309 431 633 990 608 53 146 705 889 786 888 717 441 822 43 949 736 532 767 89 69 991 806 821 270 823 793 704 621 21 658 992 137 855 291 907 788 880 506 562 59 432 475 560 773 4 105 619 329 476 228 862 558 565 830 776 628 236 256 309 755 247 757 394 554 812 198 749 731 119 561 797 10 447 856 343 843 954 672 692 131 400 638 276 660 124 393 81 829 601 339 941 188 88 515 351 191 175 514 610 146 100 164 736 846 545 336 448 711 877 403 99 554 747 266 96 325 609 34 882 876 760 728 940 810 644 865 857 368 616 257 768 595 18 295 102 657 844 774 640 796 736 9 704 365 116 970 521 209 521 788 401 770 929 726 42 702 159 830 521 551 906 353 527 996 551 836 422 714 284 105 878 855 594 467 88 507 830 747 493 32 905 819 289 187 277 749 1 652 687 880 646 254 937 153 60 815 327 424 917 752 47 398 370 905 890 249 136 185 412 905 427 974 267 305 340 736 946 227 977 488 916 297 802 321 23 103 978 900 93 132 742 923 540 502 778 253 892 227 645 471 120 209 279 358 439 562 787 576 170 875 473 207 845 224 123 605 312 142 175 223 580 315 855 554 486 125 234 208 828 488 1 367 742 418 347 222 26 269 37 243 787 65 668 952 883 786 224 726 229 865 157 830 490 832 651 347 230 215 916 932 940 680 451 6 36 401 301 359 310 926 656 33 156 291 899 549 266 372 171 423 488 498 622 788 469 689 481 337 678 429 236 623 25 223 32 487 912 521 88 952 183 822 782 783 364 507 598 260 294 34 413 607 801 271 3 190 72 815 649 207 484 987 64 454 765 581 678 330 399 733 366 826 753 895 383 922 325 890 601 760 980 761 767 555 420 148 601 204 448 431 54 581 616 261 196 325 248 511 576 692 385 399 781 551 814 154 636 758 343 603 700 875 935 327 494 450 44 181 717 121 487 551 487 295 210 85 591 584 847 956 98 903 458 843 403 983 652 899 830 896 41 775 933 798 78 168 858 670 309 600 966 527 992 149 667 680 82 285 639 949 305 768 306 72 455 918 92 281 196 964 977 603 624 694 982 687 259 910 722 413 9 874 663 926 962 810 916 456 369 74 502 310 803 827 693 941 963 992 894 609 302 470 957 758 819 902 629 306 351 387 478 326 946 135 58 963 49 496 145 301 614 48 568 103 899 82 819 756 148 96 496 866 911 942 817 994 368 143 379 530 229 100 273 991 251 370 233 278 685 573 81 998 66 33 239 224 930 779 396 105 535 737 370 606 399 937 511 789 393 11 949 654 376 1 13 521 182 18 780 211 246 871 920 452 992 637 792 263 183 117 485 62 929 837 124 482 148 736 961 739 354 174 896 694 151 73 992 560 407 490 804 699 324 917 991 380 154 89 89 460 320 599 40 787 274 505 384 590 474 843 969 625 100 692 958 541 527 756 780 102 35 354 352 861 171 194 616 397 77 989 425 72 856 129 957 130 24 935 7 999 6 549 472 219 2 833 532 708 173 730 27 55 238 60 524 185 929 441 80 964 613 687 778 996 93 946 778 432 687 33 503 42 753 70 365 577 257 254 709 374 725 290 451 128 870 409 437 828 370 632 149 751 202 521 734 99 882 231 118 970 439 995 403 850 829 275 18 21 975 573 553 997 199 618 459 899 796 911 433 183 255 266 103 475 837 270 898 17 857 612 103 688 944 460 682 466 781 461 461 877 224 423 919 575 610 950 986 9 411 537 257 885 179 305 428 316 378 617 994 952 305 835 433 346 43 438 866 382 532 758 277 618 941 954 503 524 712 728 465 592 17 651 964 667 961 370 234 46 783 802 235 319 367 276 146 842 74 621 837 241 858 545 115 523 289 196 180 64 106 248 232 783 407 513 552 735 224 641 137 446 9 175 119 31 580 989 498 786 540 648 733 656 452 917 254 759 112 647 831 941 620 874 580 309 948 741 840 185 672 228 689 558 367